// vim: sw=4 ts=4 et
// Eagle scaler
//
// This implements Eagle, as described by Dirk Stevens, as well as Scale2x.
//
// Basic operation:
//
//   Eagle and Scale2x are both doubling algorithms working pixel-by-pixel.  They operate on a
//   matrix as such:
//
//      -1 0 1 2
//  -1   I E F J
//   0   G A B K  =>  A'  A'''
//   1   H C D L      A'' A''''
//   2   M N O P
//
// Eagle:
//
//  I E F    A'   A'''    A'  <= G==I==E ? I : A     A'''  <= E==F==B ? F : A
//  G A B => A''  A''''   A'' <= C==H==G ? H : A     A'''' <= B==D==C ? Z : A
//  H C D
//
//  Pathology:  if all but A are the same color, A vanishes.
//
// Scale2x:
//
//    E        A'   A'''
//  G A B  =>  A''  A''''
//    C
//
//  Match[1] <= G==E    A'    <= Match[1] ? E : A
//  Match[2] <= E==B    A''   <= Match[2] ? B : A
//  Match[3] <= B==C    A'''  <= Match[3] ? C : A
//  Match[4] <= C==G    A'''' <= Match[4] ? G : A
//
//  If fewer than two mismatch, set all 4 to A.  Avoids Eagle pathology:
//  if ( !(
//       (!Match[1] && !(Match[2] && Match[3] && Match[4]))
//    || (!Match[2] && !(Match[3] && Match[4]))
//    || (!Match[3] && !Match[4]))
//        )
//   A' <= A; A'' <= A; A''' <= A; A'''' <= A
//
// Scale3x:
//
//  I E F    A'1  A'4  A'7
//  G A B => A'2  A    A'8
//  H C D    A'3  A'6  A'9
//
// Observations:
//  - Eagle adds the corner to Scale2x Match[n] and, if matching, selects the corner
//  - Scale2x pathology avoidance can be applied to Eagle
//  - Scale2x uses the corner for calculations, but selects from the sides
//  - All output pixels are generated by relationships not easily replicated by muxes, so the least
//    logic and routing is used by computing all outputs on the same clock in parallel
//  - Expanding one pixel requires 27 bytes for 24-bit color input, plus 27 bytes for 3x3 output;
//    managing this from a BRAM is hard, but 3 lines of 1920 at 24 bits is over 16KiB.  For 2xSaI,
//    it approaches 30KiB including transparency.  This block RAM should be shared for use by the
//    selected filter, and must be divided up to allow 96 bits (12 bytes) access simultaneously on
//    each clock so as to rotate the input filter.