// vim: sw=4 ts=4 et
// Interfaces to the ASCAL Avalon Scaler
//
// License: MIT